//-----------------------------------------------------------------------
//	File:		$RCSfile: VideoROM.v,v $
//	Version:	$Revision: 1.2 $
//	Desc:		ITU656/601 Video Test ROM
//	Author:		Greg Gibeling
//	Copyright:	Copyright 2003 UC Berkeley
//	This copyright header must appear in all derivative works.
//-----------------------------------------------------------------------

//-----------------------------------------------------------------------
//	Section:	Change Log
//-----------------------------------------------------------------------
//	$Log: VideoROM.v,v $
//	Revision 1.2  2004/10/05 20:00:16  Administrator
//	Fixed module name bug
//	
//	Revision 1.1  2004/10/05 19:56:01  SYSTEM
//	Initial Import
//	
//-----------------------------------------------------------------------

//-----------------------------------------------------------------------
//	Section:	Includes
//-----------------------------------------------------------------------
`include "Const.v"
//-----------------------------------------------------------------------

//-----------------------------------------------------------------------
//	Module:		VideoROM
//	Desc:		This module generates a series of solid color
//			bars as a test pattern.
//	Params:		totallines:	The total number of video lines
//					to output.
//			activelines:	The total number of active video
//					lines to output
//			f0topblank:	The number of vertical blanking
//					lines to insert above the active
//					portion of the 0 (Odd) field.
//			hblanksamples:	The number of samples (16bit
//					words) per line which are
//					blanking.  Includes SAV/EAV
//			activesamples:	The number of active video samples
//					per line.
//-----------------------------------------------------------------------
module	VideoROM(	//-----------------------------------------------
			//	System Inputs
			//-----------------------------------------------
			Clock,
			Reset,
			//-----------------------------------------------

			//-----------------------------------------------
			//	Video Data Host Interface
			//-----------------------------------------------
			DOut,
			OutRequest,
			OutRequestLine,
			OutRequestPair
			//-----------------------------------------------
		);


	//---------------------------------------------------------------
	//	System Inputs
	//---------------------------------------------------------------
	input			Clock, Reset;
	//---------------------------------------------------------------

	//---------------------------------------------------------------
	//	Video Data Host Interface
	//---------------------------------------------------------------
	output	[31:0]		DOut;
	input			OutRequest;
	input	[8:0]	OutRequestLine;
	input	[8:0]	OutRequestPair;
	//---------------------------------------------------------------

	//---------------------------------------------------------------
	//	Regs
	//---------------------------------------------------------------
	reg	[31:0]		DOutRaw;
	reg					Pipe;
	
	always @ (posedge Clock) begin
		if(Reset)
			Pipe <= 1'b0;
		else if(OutRequest)
			Pipe <= 1'b1;
		else
			Pipe <= 1'b0;
	
	end
	
	//---------------------------------------------------------------
	//	Test Video Generator
	//---------------------------------------------------------------
	always @ ( * ) begin
		DOutRaw = 32'h10801080;
		
		if((OutRequestLine >> 2) == 6) begin
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 51)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 53)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 54)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 55)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 56)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 79)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 80)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 81)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 84)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 88)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 93)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 95)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 97)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 106)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 7) begin
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 56)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 84)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 8) begin
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 56)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 84)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 9) begin
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 57)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 84)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 10) begin
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 57)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 79)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 80)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 81)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 84)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 88)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 97)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 11) begin
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 57)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 12) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 58)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 13) begin
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 53)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 58)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 14) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 53)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 58)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 15) begin
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 53)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 59)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 16) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 53)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 54)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 59)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 17) begin
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 59)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 18) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 60)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 19) begin
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 60)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 20) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 60)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 111)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 112)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 114)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 121)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 21) begin
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 22) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 51)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 53)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 54)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 55)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 56)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 23) begin
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 56)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 24) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 57)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 58)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 59)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 60)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 93)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 95)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 106)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 111)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 112)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 114)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 121)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 25) begin
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 26) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 27) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 28) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 79)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 80)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 81)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 83)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 84)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 88)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 111)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 112)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 114)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 121)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 29) begin
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 143)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 30) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 143)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 144)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 31) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 144)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 32) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 79)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 80)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 81)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 83)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 84)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 111)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 112)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 121)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 145)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 33) begin
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 145)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 34) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 145)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 35) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 93)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 95)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 97)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 145)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 36) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 79)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 144)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 37) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 80)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 81)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 143)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 144)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 38) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 83)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 143)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 39) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 84)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 93)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 95)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 97)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 40) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 41) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 42) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 79)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 111)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 112)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 121)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 43) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 44) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 84)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 45) begin
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 83)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 84)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 46) begin
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 79)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 80)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 81)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 88)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 111)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 112)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 114)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 121)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 47) begin
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 51)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 53)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 54)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 55)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 48) begin
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 51)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 53)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 54)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 55)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 56)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 49) begin
			if(OutRequestPair>>1 == 51)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 53)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 54)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 55)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 56)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 57)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 58)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 59)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 50) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 54)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 55)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 56)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 57)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 58)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 59)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 60)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 51) begin
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 56)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 57)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 58)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 59)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 60)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 52) begin
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 57)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 58)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 59)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 60)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 53) begin
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 59)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 60)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h15801580;
		end

		if((OutRequestLine >> 2) == 54) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 60)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 55) begin
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 56) begin
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 57) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h15801580;
		end

		if((OutRequestLine >> 2) == 58) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 59) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 60) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 61) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 62) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 51)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 63) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 51)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 64) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 51)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 65) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 51)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 66) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 67) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 68) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 52)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 69) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 70) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 71) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 72) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 73) begin
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 74) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 75) begin
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 76) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 77) begin
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 78) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 79) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 80) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 60)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 81) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 59)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 82) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 58)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 60)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 83) begin
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 59)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 84) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 58)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 60)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 85) begin
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 57)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 88)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 93)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 106)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 111)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 112)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 114)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 86) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 61)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 95)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 87) begin
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 88) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 40)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 41)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 42)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 43)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 44)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 50)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 62)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 63)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 93)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 114)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 89) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 45)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 46)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 47)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 106)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 90) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 64)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 77)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 93)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 114)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 91) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 48)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 49)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 65)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 79)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 95)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 92) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'h758b7580;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 66)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 68)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 70)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 78)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 79)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 93)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 106)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 114)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 93) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 67)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 69)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 71)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 79)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 94) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 72)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 79)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 80)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 106)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 114)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 95) begin
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'h758b7580;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 73)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 79)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 131)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 96) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 12)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h758b7580;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 74)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 75)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 76)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 80)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 88)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 106)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 107)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 111)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 112)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 114)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 119)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 97) begin
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 13)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 80)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 81)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 98) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 16)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'h758b7580;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 80)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 81)
				DOutRaw = 32'h2f802f92;
		end

		if((OutRequestLine >> 2) == 99) begin
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 11)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 17)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 18)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 19)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 20)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 21)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 81)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 88)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 93)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 97)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 106)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 112)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 114)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 121)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 100) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 10)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 14)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 15)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 22)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 81)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 106)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 111)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 101) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 23)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 81)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 106)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 111)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 102) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 8)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 24)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'h758b7580;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 93)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 96)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 97)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 98)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 104)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 105)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 106)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 132)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 133)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 134)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 140)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 141)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 142)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 103) begin
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 7)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 9)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 104) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h40854080;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 6)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 25)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 82)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 105) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 5)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 83)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 93)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 112)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 106) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 26)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h758b7580;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 83)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 88)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 107) begin
			if(OutRequestPair>>1 == 27)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 29)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'h758b7580;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 83)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 95)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 108) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 28)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 30)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h758b7580;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h758b7580;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 84)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 88)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 95)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 124)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 109) begin
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'h758b7580;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 95)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 111)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 112)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 113)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 114)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 125)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 110) begin
			if(OutRequestPair>>1 == 4)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 31)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'hb080b0d3;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 84)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 86)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 87)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 88)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 89)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 90)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 91)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 92)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 93)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 94)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 99)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 100)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 101)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 102)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 103)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 108)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 109)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 110)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 111)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 115)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 116)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 117)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 118)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 120)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 121)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 122)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 123)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 126)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 127)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 128)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 129)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 130)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 135)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 136)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 137)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 138)
				DOutRaw = 32'hcd96cd80;
			if(OutRequestPair>>1 == 139)
				DOutRaw = 32'hcd96cd80;
		end

		if((OutRequestLine >> 2) == 111) begin
			if(OutRequestPair>>1 == 32)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 33)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 34)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 35)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 36)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 37)
				DOutRaw = 32'h5f805fb0;
			if(OutRequestPair>>1 == 38)
				DOutRaw = 32'h15801580;
			if(OutRequestPair>>1 == 39)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 83)
				DOutRaw = 32'h2f802f92;
			if(OutRequestPair>>1 == 85)
				DOutRaw = 32'h2f802f92;
		end


	end
	//---------------------------------------------------------------

	//---------------------------------------------------------------
	//	Output Register
	//---------------------------------------------------------------
	Register	DOReg(	.Clock(		Clock),
				.Reset(		Reset),
				.Set(		1'b0),
				.Enable(	Pipe),
				.In(		DOutRaw),
				.Out(		DOut));
	defparam	DOReg.width =		32;
	//---------------------------------------------------------------
endmodule
//-----------------------------------------------------------------------