module PlaceWriteFSM(Clock, Reset, WEn, Length, WRow, WCol);

endmodule